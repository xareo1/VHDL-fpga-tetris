library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package AUDIO_PACKAGE is

    constant NOTE_COUNT : INTEGER := 384;
    type ROM_AUDIO is array (0 to 383) of INTEGER;
    
    constant pitch_rom : ROM_AUDIO :=
    (
        0 => 75872 - 1,
        1 => 303030 - 1,
        2 => 101214 - 1,
        3 => 95602 - 1,
        4 => 85178 - 1,
        5 => 75872 - 1,
        6 => 85178 - 1,
        7 => 95602 - 1,
        8 => 101214 - 1,
        9 => 113636 - 1,
        10 => 227272 - 1,
        11 => 113636 - 1,
        12 => 95602 - 1,
        13 => 75872 - 1,
        14 => 227272 - 1,
        15 => 85178 - 1,
        16 => 95602 - 1,
        17 => 101214 - 1,
        18 => 151515 - 1,
        19 => 127551 - 1,
        20 => 95602 - 1,
        21 => 85178 - 1,
        22 => 303030 - 1,
        23 => 75872 - 1,
        24 => 303030 - 1,
        25 => 95602 - 1,
        26 => 227272 - 1,
        27 => 113636 - 1,
        28 => 227272 - 1,
        29 => 113636 - 1,
        30 => 227272 - 1,
        31 => 406504 - 1,
        32 => 381679 - 1,
        33 => 340136 - 1,
        34 => 85178 - 1,
        35 => 71633 - 1,
        36 => 56818 - 1,
        37 => 95602 - 1,
        38 => 95602 - 1,
        39 => 63775 - 1,
        40 => 71633 - 1,
        41 => 75872 - 1,
        42 => 381679 - 1,
        43 => 100000000 - 1,
        44 => 95602 - 1,
        45 => 75872 - 1,
        46 => 113636 - 1,
        47 => 127551 - 1,
        48 => 85178 - 1,
        49 => 95602 - 1,
        50 => 101214 - 1,
        51 => 151515 - 1,
        52 => 101214 - 1,
        53 => 95602 - 1,
        54 => 85178 - 1,
        55 => 127551 - 1,
        56 => 75872 - 1,
        57 => 127551 - 1,
        58 => 95602 - 1,
        59 => 151515 - 1,
        60 => 113636 - 1,
        61 => 303030 - 1,
        62 => 113636 - 1,
        63 => 100000000 - 1,
        64 => 75872 - 1,
        65 => 303030 - 1,
        66 => 101214 - 1,
        67 => 95602 - 1,
        68 => 85178 - 1,
        69 => 75872 - 1,
        70 => 85178 - 1,
        71 => 95602 - 1,
        72 => 101214 - 1,
        73 => 113636 - 1,
        74 => 227272 - 1,
        75 => 113636 - 1,
        76 => 95602 - 1,
        77 => 75872 - 1,
        78 => 227272 - 1,
        79 => 85178 - 1,
        80 => 95602 - 1,
        81 => 101214 - 1,
        82 => 151515 - 1,
        83 => 127551 - 1,
        84 => 95602 - 1,
        85 => 85178 - 1,
        86 => 303030 - 1,
        87 => 75872 - 1,
        88 => 303030 - 1,
        89 => 95602 - 1,
        90 => 227272 - 1,
        91 => 113636 - 1,
        92 => 227272 - 1,
        93 => 113636 - 1,
        94 => 227272 - 1,
        95 => 406504 - 1,
        96 => 381679 - 1,
        97 => 340136 - 1,
        98 => 85178 - 1,
        99 => 71633 - 1,
        100 => 56818 - 1,
        101 => 95602 - 1,
        102 => 95602 - 1,
        103 => 63775 - 1,
        104 => 71633 - 1,
        105 => 75872 - 1,
        106 => 381679 - 1,
        107 => 100000000 - 1,
        108 => 95602 - 1,
        109 => 75872 - 1,
        110 => 113636 - 1,
        111 => 127551 - 1,
        112 => 85178 - 1,
        113 => 95602 - 1,
        114 => 101214 - 1,
        115 => 151515 - 1,
        116 => 101214 - 1,
        117 => 95602 - 1,
        118 => 85178 - 1,
        119 => 127551 - 1,
        120 => 75872 - 1,
        121 => 127551 - 1,
        122 => 95602 - 1,
        123 => 151515 - 1,
        124 => 113636 - 1,
        125 => 303030 - 1,
        126 => 113636 - 1,
        127 => 100000000 - 1,
        128 => 151515 - 1,
        129 => 303030 - 1,
        130 => 454545 - 1,
        131 => 303030 - 1,
        132 => 190839 - 1,
        133 => 303030 - 1,
        134 => 454545 - 1,
        135 => 303030 - 1,
        136 => 170068 - 1,
        137 => 303030 - 1,
        138 => 480769 - 1,
        139 => 303030 - 1,
        140 => 202429 - 1,
        141 => 303030 - 1,
        142 => 480769 - 1,
        143 => 303030 - 1,
        144 => 190839 - 1,
        145 => 303030 - 1,
        146 => 454545 - 1,
        147 => 303030 - 1,
        148 => 227272 - 1,
        149 => 303030 - 1,
        150 => 454545 - 1,
        151 => 303030 - 1,
        152 => 240384 - 1,
        153 => 303030 - 1,
        154 => 480769 - 1,
        155 => 303030 - 1,
        156 => 202429 - 1,
        157 => 303030 - 1,
        158 => 480769 - 1,
        159 => 303030 - 1,
        160 => 151515 - 1,
        161 => 303030 - 1,
        162 => 454545 - 1,
        163 => 303030 - 1,
        164 => 190839 - 1,
        165 => 303030 - 1,
        166 => 454545 - 1,
        167 => 303030 - 1,
        168 => 170068 - 1,
        169 => 303030 - 1,
        170 => 480769 - 1,
        171 => 303030 - 1,
        172 => 202429 - 1,
        173 => 303030 - 1,
        174 => 480769 - 1,
        175 => 303030 - 1,
        176 => 190839 - 1,
        177 => 303030 - 1,
        178 => 151515 - 1,
        179 => 303030 - 1,
        180 => 113636 - 1,
        181 => 303030 - 1,
        182 => 454545 - 1,
        183 => 303030 - 1,
        184 => 120481 - 1,
        185 => 303030 - 1,
        186 => 480769 - 1,
        187 => 303030 - 1,
        188 => 480769 - 1,
        189 => 303030 - 1,
        190 => 480769 - 1,
        191 => 303030 - 1,
        192 => 75872 - 1,
        193 => 303030 - 1,
        194 => 101214 - 1,
        195 => 95602 - 1,
        196 => 85178 - 1,
        197 => 75872 - 1,
        198 => 85178 - 1,
        199 => 95602 - 1,
        200 => 101214 - 1,
        201 => 113636 - 1,
        202 => 227272 - 1,
        203 => 113636 - 1,
        204 => 95602 - 1,
        205 => 75872 - 1,
        206 => 227272 - 1,
        207 => 85178 - 1,
        208 => 95602 - 1,
        209 => 101214 - 1,
        210 => 151515 - 1,
        211 => 127551 - 1,
        212 => 95602 - 1,
        213 => 85178 - 1,
        214 => 303030 - 1,
        215 => 75872 - 1,
        216 => 303030 - 1,
        217 => 95602 - 1,
        218 => 227272 - 1,
        219 => 113636 - 1,
        220 => 227272 - 1,
        221 => 113636 - 1,
        222 => 227272 - 1,
        223 => 406504 - 1,
        224 => 381679 - 1,
        225 => 340136 - 1,
        226 => 85178 - 1,
        227 => 71633 - 1,
        228 => 56818 - 1,
        229 => 95602 - 1,
        230 => 95602 - 1,
        231 => 63775 - 1,
        232 => 71633 - 1,
        233 => 75872 - 1,
        234 => 381679 - 1,
        235 => 100000000 - 1,
        236 => 95602 - 1,
        237 => 75872 - 1,
        238 => 113636 - 1,
        239 => 127551 - 1,
        240 => 85178 - 1,
        241 => 95602 - 1,
        242 => 101214 - 1,
        243 => 151515 - 1,
        244 => 101214 - 1,
        245 => 95602 - 1,
        246 => 85178 - 1,
        247 => 127551 - 1,
        248 => 75872 - 1,
        249 => 127551 - 1,
        250 => 95602 - 1,
        251 => 151515 - 1,
        252 => 113636 - 1,
        253 => 303030 - 1,
        254 => 113636 - 1,
        255 => 100000000 - 1,
        256 => 75872 - 1,
        257 => 303030 - 1,
        258 => 101214 - 1,
        259 => 95602 - 1,
        260 => 85178 - 1,
        261 => 75872 - 1,
        262 => 85178 - 1,
        263 => 95602 - 1,
        264 => 101214 - 1,
        265 => 113636 - 1,
        266 => 227272 - 1,
        267 => 113636 - 1,
        268 => 95602 - 1,
        269 => 75872 - 1,
        270 => 227272 - 1,
        271 => 85178 - 1,
        272 => 95602 - 1,
        273 => 101214 - 1,
        274 => 151515 - 1,
        275 => 127551 - 1,
        276 => 95602 - 1,
        277 => 85178 - 1,
        278 => 303030 - 1,
        279 => 75872 - 1,
        280 => 303030 - 1,
        281 => 95602 - 1,
        282 => 227272 - 1,
        283 => 113636 - 1,
        284 => 227272 - 1,
        285 => 113636 - 1,
        286 => 227272 - 1,
        287 => 406504 - 1,
        288 => 381679 - 1,
        289 => 340136 - 1,
        290 => 85178 - 1,
        291 => 71633 - 1,
        292 => 56818 - 1,
        293 => 95602 - 1,
        294 => 95602 - 1,
        295 => 63775 - 1,
        296 => 71633 - 1,
        297 => 75872 - 1,
        298 => 381679 - 1,
        299 => 100000000 - 1,
        300 => 95602 - 1,
        301 => 75872 - 1,
        302 => 113636 - 1,
        303 => 127551 - 1,
        304 => 85178 - 1,
        305 => 95602 - 1,
        306 => 101214 - 1,
        307 => 151515 - 1,
        308 => 101214 - 1,
        309 => 95602 - 1,
        310 => 85178 - 1,
        311 => 127551 - 1,
        312 => 75872 - 1,
        313 => 127551 - 1,
        314 => 95602 - 1,
        315 => 151515 - 1,
        316 => 113636 - 1,
        317 => 303030 - 1,
        318 => 113636 - 1,
        319 => 100000000 - 1,
        320 => 151515 - 1,
        321 => 303030 - 1,
        322 => 454545 - 1,
        323 => 303030 - 1,
        324 => 190839 - 1,
        325 => 303030 - 1,
        326 => 454545 - 1,
        327 => 303030 - 1,
        328 => 170068 - 1,
        329 => 303030 - 1,
        330 => 480769 - 1,
        331 => 303030 - 1,
        332 => 202429 - 1,
        333 => 303030 - 1,
        334 => 480769 - 1,
        335 => 303030 - 1,
        336 => 190839 - 1,
        337 => 303030 - 1,
        338 => 454545 - 1,
        339 => 303030 - 1,
        340 => 227272 - 1,
        341 => 303030 - 1,
        342 => 454545 - 1,
        343 => 303030 - 1,
        344 => 240384 - 1,
        345 => 303030 - 1,
        346 => 480769 - 1,
        347 => 303030 - 1,
        348 => 202429 - 1,
        349 => 303030 - 1,
        350 => 480769 - 1,
        351 => 303030 - 1,
        352 => 151515 - 1,
        353 => 303030 - 1,
        354 => 454545 - 1,
        355 => 303030 - 1,
        356 => 190839 - 1,
        357 => 303030 - 1,
        358 => 454545 - 1,
        359 => 303030 - 1,
        360 => 170068 - 1,
        361 => 303030 - 1,
        362 => 480769 - 1,
        363 => 303030 - 1,
        364 => 202429 - 1,
        365 => 303030 - 1,
        366 => 480769 - 1,
        367 => 303030 - 1,
        368 => 190839 - 1,
        369 => 303030 - 1,
        370 => 151515 - 1,
        371 => 303030 - 1,
        372 => 113636 - 1,
        373 => 303030 - 1,
        374 => 454545 - 1,
        375 => 303030 - 1,
        376 => 120481 - 1,
        377 => 303030 - 1,
        378 => 480769 - 1,
        379 => 303030 - 1,
        380 => 480769 - 1,
        381 => 303030 - 1,
        382 => 480769 - 1,
        383 => 303030 - 1
    );
    
    constant duration_rom : ROM_AUDIO :=
    (
        0 => 20000000 - 1,
        1 => 20000000 - 1,
        2 => 20000000 - 1,
        3 => 20000000 - 1,
        4 => 20000000 - 1,
        5 => 10000000 - 1,
        6 => 10000000 - 1,
        7 => 20000000 - 1,
        8 => 20000000 - 1,
        9 => 20000000 - 1,
        10 => 20000000 - 1,
        11 => 20000000 - 1,
        12 => 20000000 - 1,
        13 => 20000000 - 1,
        14 => 20000000 - 1,
        15 => 20000000 - 1,
        16 => 20000000 - 1,
        17 => 20000000 - 1,
        18 => 20000000 - 1,
        19 => 20000000 - 1,
        20 => 20000000 - 1,
        21 => 20000000 - 1,
        22 => 20000000 - 1,
        23 => 20000000 - 1,
        24 => 20000000 - 1,
        25 => 20000000 - 1,
        26 => 20000000 - 1,
        27 => 20000000 - 1,
        28 => 20000000 - 1,
        29 => 20000000 - 1,
        30 => 20000000 - 1,
        31 => 20000000 - 1,
        32 => 20000000 - 1,
        33 => 20000000 - 1,
        34 => 40000000 - 1,
        35 => 20000000 - 1,
        36 => 20000000 - 1,
        37 => 10000000 - 1,
        38 => 10000000 - 1,
        39 => 20000000 - 1,
        40 => 20000000 - 1,
        41 => 20000000 - 1,
        42 => 20000000 - 1,
        43 => 20000000 - 1,
        44 => 20000000 - 1,
        45 => 20000000 - 1,
        46 => 10000000 - 1,
        47 => 10000000 - 1,
        48 => 20000000 - 1,
        49 => 20000000 - 1,
        50 => 20000000 - 1,
        51 => 20000000 - 1,
        52 => 20000000 - 1,
        53 => 20000000 - 1,
        54 => 20000000 - 1,
        55 => 20000000 - 1,
        56 => 20000000 - 1,
        57 => 20000000 - 1,
        58 => 20000000 - 1,
        59 => 20000000 - 1,
        60 => 20000000 - 1,
        61 => 20000000 - 1,
        62 => 40000000 - 1,
        63 => 40000000 - 1,
        64 => 20000000 - 1,
        65 => 20000000 - 1,
        66 => 20000000 - 1,
        67 => 20000000 - 1,
        68 => 20000000 - 1,
        69 => 10000000 - 1,
        70 => 10000000 - 1,
        71 => 20000000 - 1,
        72 => 20000000 - 1,
        73 => 20000000 - 1,
        74 => 20000000 - 1,
        75 => 20000000 - 1,
        76 => 20000000 - 1,
        77 => 20000000 - 1,
        78 => 20000000 - 1,
        79 => 20000000 - 1,
        80 => 20000000 - 1,
        81 => 20000000 - 1,
        82 => 20000000 - 1,
        83 => 20000000 - 1,
        84 => 20000000 - 1,
        85 => 20000000 - 1,
        86 => 20000000 - 1,
        87 => 20000000 - 1,
        88 => 20000000 - 1,
        89 => 20000000 - 1,
        90 => 20000000 - 1,
        91 => 20000000 - 1,
        92 => 20000000 - 1,
        93 => 20000000 - 1,
        94 => 20000000 - 1,
        95 => 20000000 - 1,
        96 => 20000000 - 1,
        97 => 20000000 - 1,
        98 => 40000000 - 1,
        99 => 20000000 - 1,
        100 => 20000000 - 1,
        101 => 10000000 - 1,
        102 => 10000000 - 1,
        103 => 20000000 - 1,
        104 => 20000000 - 1,
        105 => 20000000 - 1,
        106 => 20000000 - 1,
        107 => 20000000 - 1,
        108 => 20000000 - 1,
        109 => 20000000 - 1,
        110 => 10000000 - 1,
        111 => 10000000 - 1,
        112 => 20000000 - 1,
        113 => 20000000 - 1,
        114 => 20000000 - 1,
        115 => 20000000 - 1,
        116 => 20000000 - 1,
        117 => 20000000 - 1,
        118 => 20000000 - 1,
        119 => 20000000 - 1,
        120 => 20000000 - 1,
        121 => 20000000 - 1,
        122 => 20000000 - 1,
        123 => 20000000 - 1,
        124 => 20000000 - 1,
        125 => 20000000 - 1,
        126 => 40000000 - 1,
        127 => 40000000 - 1,
        128 => 20000000 - 1,
        129 => 20000000 - 1,
        130 => 20000000 - 1,
        131 => 20000000 - 1,
        132 => 20000000 - 1,
        133 => 20000000 - 1,
        134 => 20000000 - 1,
        135 => 20000000 - 1,
        136 => 20000000 - 1,
        137 => 20000000 - 1,
        138 => 20000000 - 1,
        139 => 20000000 - 1,
        140 => 20000000 - 1,
        141 => 20000000 - 1,
        142 => 20000000 - 1,
        143 => 20000000 - 1,
        144 => 20000000 - 1,
        145 => 20000000 - 1,
        146 => 20000000 - 1,
        147 => 20000000 - 1,
        148 => 20000000 - 1,
        149 => 20000000 - 1,
        150 => 20000000 - 1,
        151 => 20000000 - 1,
        152 => 20000000 - 1,
        153 => 20000000 - 1,
        154 => 20000000 - 1,
        155 => 20000000 - 1,
        156 => 20000000 - 1,
        157 => 20000000 - 1,
        158 => 20000000 - 1,
        159 => 20000000 - 1,
        160 => 20000000 - 1,
        161 => 20000000 - 1,
        162 => 20000000 - 1,
        163 => 20000000 - 1,
        164 => 20000000 - 1,
        165 => 20000000 - 1,
        166 => 20000000 - 1,
        167 => 20000000 - 1,
        168 => 20000000 - 1,
        169 => 20000000 - 1,
        170 => 20000000 - 1,
        171 => 20000000 - 1,
        172 => 20000000 - 1,
        173 => 20000000 - 1,
        174 => 20000000 - 1,
        175 => 20000000 - 1,
        176 => 20000000 - 1,
        177 => 20000000 - 1,
        178 => 20000000 - 1,
        179 => 20000000 - 1,
        180 => 20000000 - 1,
        181 => 20000000 - 1,
        182 => 20000000 - 1,
        183 => 20000000 - 1,
        184 => 20000000 - 1,
        185 => 20000000 - 1,
        186 => 20000000 - 1,
        187 => 20000000 - 1,
        188 => 20000000 - 1,
        189 => 20000000 - 1,
        190 => 20000000 - 1,
        191 => 20000000 - 1,
        192 => 20000000 - 1,
        193 => 20000000 - 1,
        194 => 20000000 - 1,
        195 => 20000000 - 1,
        196 => 20000000 - 1,
        197 => 10000000 - 1,
        198 => 10000000 - 1,
        199 => 20000000 - 1,
        200 => 20000000 - 1,
        201 => 20000000 - 1,
        202 => 20000000 - 1,
        203 => 20000000 - 1,
        204 => 20000000 - 1,
        205 => 20000000 - 1,
        206 => 20000000 - 1,
        207 => 20000000 - 1,
        208 => 20000000 - 1,
        209 => 20000000 - 1,
        210 => 20000000 - 1,
        211 => 20000000 - 1,
        212 => 20000000 - 1,
        213 => 20000000 - 1,
        214 => 20000000 - 1,
        215 => 20000000 - 1,
        216 => 20000000 - 1,
        217 => 20000000 - 1,
        218 => 20000000 - 1,
        219 => 20000000 - 1,
        220 => 20000000 - 1,
        221 => 20000000 - 1,
        222 => 20000000 - 1,
        223 => 20000000 - 1,
        224 => 20000000 - 1,
        225 => 20000000 - 1,
        226 => 40000000 - 1,
        227 => 20000000 - 1,
        228 => 20000000 - 1,
        229 => 10000000 - 1,
        230 => 10000000 - 1,
        231 => 20000000 - 1,
        232 => 20000000 - 1,
        233 => 20000000 - 1,
        234 => 20000000 - 1,
        235 => 20000000 - 1,
        236 => 20000000 - 1,
        237 => 20000000 - 1,
        238 => 10000000 - 1,
        239 => 10000000 - 1,
        240 => 20000000 - 1,
        241 => 20000000 - 1,
        242 => 20000000 - 1,
        243 => 20000000 - 1,
        244 => 20000000 - 1,
        245 => 20000000 - 1,
        246 => 20000000 - 1,
        247 => 20000000 - 1,
        248 => 20000000 - 1,
        249 => 20000000 - 1,
        250 => 20000000 - 1,
        251 => 20000000 - 1,
        252 => 20000000 - 1,
        253 => 20000000 - 1,
        254 => 40000000 - 1,
        255 => 40000000 - 1,
        256 => 20000000 - 1,
        257 => 20000000 - 1,
        258 => 20000000 - 1,
        259 => 20000000 - 1,
        260 => 20000000 - 1,
        261 => 10000000 - 1,
        262 => 10000000 - 1,
        263 => 20000000 - 1,
        264 => 20000000 - 1,
        265 => 20000000 - 1,
        266 => 20000000 - 1,
        267 => 20000000 - 1,
        268 => 20000000 - 1,
        269 => 20000000 - 1,
        270 => 20000000 - 1,
        271 => 20000000 - 1,
        272 => 20000000 - 1,
        273 => 20000000 - 1,
        274 => 20000000 - 1,
        275 => 20000000 - 1,
        276 => 20000000 - 1,
        277 => 20000000 - 1,
        278 => 20000000 - 1,
        279 => 20000000 - 1,
        280 => 20000000 - 1,
        281 => 20000000 - 1,
        282 => 20000000 - 1,
        283 => 20000000 - 1,
        284 => 20000000 - 1,
        285 => 20000000 - 1,
        286 => 20000000 - 1,
        287 => 20000000 - 1,
        288 => 20000000 - 1,
        289 => 20000000 - 1,
        290 => 40000000 - 1,
        291 => 20000000 - 1,
        292 => 20000000 - 1,
        293 => 10000000 - 1,
        294 => 10000000 - 1,
        295 => 20000000 - 1,
        296 => 20000000 - 1,
        297 => 20000000 - 1,
        298 => 20000000 - 1,
        299 => 20000000 - 1,
        300 => 20000000 - 1,
        301 => 20000000 - 1,
        302 => 10000000 - 1,
        303 => 10000000 - 1,
        304 => 20000000 - 1,
        305 => 20000000 - 1,
        306 => 20000000 - 1,
        307 => 20000000 - 1,
        308 => 20000000 - 1,
        309 => 20000000 - 1,
        310 => 20000000 - 1,
        311 => 20000000 - 1,
        312 => 20000000 - 1,
        313 => 20000000 - 1,
        314 => 20000000 - 1,
        315 => 20000000 - 1,
        316 => 20000000 - 1,
        317 => 20000000 - 1,
        318 => 40000000 - 1,
        319 => 40000000 - 1,
        320 => 20000000 - 1,
        321 => 20000000 - 1,
        322 => 20000000 - 1,
        323 => 20000000 - 1,
        324 => 20000000 - 1,
        325 => 20000000 - 1,
        326 => 20000000 - 1,
        327 => 20000000 - 1,
        328 => 20000000 - 1,
        329 => 20000000 - 1,
        330 => 20000000 - 1,
        331 => 20000000 - 1,
        332 => 20000000 - 1,
        333 => 20000000 - 1,
        334 => 20000000 - 1,
        335 => 20000000 - 1,
        336 => 20000000 - 1,
        337 => 20000000 - 1,
        338 => 20000000 - 1,
        339 => 20000000 - 1,
        340 => 20000000 - 1,
        341 => 20000000 - 1,
        342 => 20000000 - 1,
        343 => 20000000 - 1,
        344 => 20000000 - 1,
        345 => 20000000 - 1,
        346 => 20000000 - 1,
        347 => 20000000 - 1,
        348 => 20000000 - 1,
        349 => 20000000 - 1,
        350 => 20000000 - 1,
        351 => 20000000 - 1,
        352 => 20000000 - 1,
        353 => 20000000 - 1,
        354 => 20000000 - 1,
        355 => 20000000 - 1,
        356 => 20000000 - 1,
        357 => 20000000 - 1,
        358 => 20000000 - 1,
        359 => 20000000 - 1,
        360 => 20000000 - 1,
        361 => 20000000 - 1,
        362 => 20000000 - 1,
        363 => 20000000 - 1,
        364 => 20000000 - 1,
        365 => 20000000 - 1,
        366 => 20000000 - 1,
        367 => 20000000 - 1,
        368 => 20000000 - 1,
        369 => 20000000 - 1,
        370 => 20000000 - 1,
        371 => 20000000 - 1,
        372 => 20000000 - 1,
        373 => 20000000 - 1,
        374 => 20000000 - 1,
        375 => 20000000 - 1,
        376 => 20000000 - 1,
        377 => 20000000 - 1,
        378 => 20000000 - 1,
        379 => 20000000 - 1,
        380 => 20000000 - 1,
        381 => 20000000 - 1,
        382 => 20000000 - 1,
        383 => 20000000 - 1
    );
    
end package;
